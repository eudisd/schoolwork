library ieee;
use ieee.std_logic_1164.all;

entity addsub is
	port();
end addsub;

architecture addsub_arch of addsub is 
begin
end addsub_arch;