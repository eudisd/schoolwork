library ieee;
use ieee.std_logic_1164.all;

entity display_mouse is
	port();
end display_mouse;


architecture arch of display_mouse is 

begin


end arch;