library ieee;
use ieee.std_logic_1164.all;

entity test_control_unit is
    port();
end test_control_unit;

architecture test_arch of test_control_unit is
begin

end test_arch;

