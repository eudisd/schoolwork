library ieee;
use ieee.std_logic_1164.all;

entity control_unit is
	port();
end control_unit;

architecture control_arch of control_unit is

begin

end contro_arch;