library ieee;
use ieee.std_logic_1164.all;

entity test_cpu is
    port();
end test_cpu;

architecture test_arch of test_cpu is
begin
end test_cpu;
