library ieee;
use ieee.std_logic_1164.all;

entity mux is
	port();
end mux;

architecture arch_mux of mux is

begin

end arch_mux;