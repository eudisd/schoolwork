library ieee;
use ieee.std_logic_1164.all;


entity cpu is
	port();
end cpu;


architecture cpu_arch of cpu is

begin

end cpu_arch;